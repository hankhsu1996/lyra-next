module m; endmodule
interface i; endinterface
program p; endprogram
