// unit error[lyra.semantic[2]]: duplicate definition `foo`
module foo; endmodule
