config my_cfg;
  design top;
endconfig
