module top;
  logic x;
  logic x;
  //    ^ error[lyra.semantic[2]]: duplicate definition
endmodule
