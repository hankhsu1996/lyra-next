module decl_test;
  wire [7:0] w;
  wire signed [15:0] s;
  logic [3:0] x, y;
  parameter DEPTH = 16;
  localparam WIDTH = 8;
endmodule
