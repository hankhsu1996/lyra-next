package r;
  typedef logic [7:0] X;
  typedef enum { X, Y } kind_t;
endpackage
