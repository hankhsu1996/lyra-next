module decl_test;
  wire [7:0] w;
  logic [3:0] x, y;
  parameter DEPTH = 16;
  localparam WIDTH = 8;
endmodule
