module b; endmodule
