module foo; endmodule
