module m;
  typedef enum { A, B, C } abc_t;
  typedef enum logic [1:0] { X, Y } xy_t;
  enum { P, Q } pq;
endmodule
