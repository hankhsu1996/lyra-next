module adder(input logic a, input logic b, output logic sum);
  assign sum = a + b;
endmodule
