// LRM 5.7.2: Real literal constants

module real_literals_test;
  real r1 = 1.2;
  real r2 = 0.1;
  real r3 = 2394.26331;
  real r4 = 1.2E12;
  real r5 = 1.30e-2;
  real r6 = 0.1e-0;
  real r7 = 23E10;
  real r8 = 29E-2;
  real r9 = 236.123_763_e-12;
endmodule
