module broken(input logic a;
  assign y = a &
endmodule
