// unit error[lyra.semantic[2]]: duplicate module
module foo; endmodule
