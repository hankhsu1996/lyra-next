module top;
  logic x, y, s;
  adder u1(.a(x), .b(y), .sum(s));
endmodule
