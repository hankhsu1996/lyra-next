package p;
  typedef enum { FALSE, TRUE } bool_t;
endpackage

package q;
  typedef enum { ORIGINAL, FALSE } teeth_t;
endpackage
