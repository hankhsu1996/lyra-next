// unit error[lyra.semantic[2]]: duplicate definition `foo`
interface foo; endinterface
