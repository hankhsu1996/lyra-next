// Package with an enum that uses range members
package my_pkg;
  typedef enum { A[2:4] } my_enum_t;
endpackage
