interface my_if;
endinterface
