program my_prog;
endprogram
