package my_pkg;
  logic [7:0] data;
  parameter WIDTH = 8;
endpackage
