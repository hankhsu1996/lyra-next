module a; endmodule
