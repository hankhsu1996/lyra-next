interface my_bus;
endinterface
