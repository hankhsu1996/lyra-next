// LRM 5.8: Time literals

module time_literals;
  realtime t1 = 2ns;
  realtime t2 = 40ps;
  realtime t3 = 1us;
  realtime t4 = 100ms;
  realtime t5 = 3s;
  realtime t6 = 10fs;
  realtime t7 = 2.1ns;
endmodule
