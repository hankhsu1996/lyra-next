module top;
  my_bus u_bus();
endmodule
