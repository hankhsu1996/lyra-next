package pkg;
  typedef bit [3:0] nibble_t;
endpackage
